module winapi
pub enum Color {
	scrollbar
	background
	activecaption
	inactivecaption
	menu
	window
	windowframe
	menutest
	windowtext
	captiontext
	activeborder
	inactiveborder
	appworkspace
	hightlight
	highlighttext
	btnface
	btnshadow
	graytext
	btntext
	inactivecaptiontext
	btnhighligh
}